--HDLRegression:TB
entity my_tb_arch is
    generic (
        GC_TESTCASE : string    := "UVVM_TB"
        );
end my_tb_arch;

